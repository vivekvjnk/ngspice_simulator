

* ---
* name: eis_control
* description: "Performs AC sweep for Electrochemical Impedance Spectroscopy (EIS)."
* input_parameters:
*   ppd: {type: int, default: 10, units: "points/decade", range: [1, 100]}
*   fmin: {type: float, default: 0.001, units: "Hz", range: [1e-6, 100.0]}
*   fmax: {type: float, default: 10000.0, units: "Hz", range: [1.0, 1e9]}
* expected_outputs:
*   - "eis_data.txt"
*   - "nyquist_plot.png"
* constraints:
*   - "fmax > fmin"
*   - "ppd > 0"
* ---




* --- control ---

* Test Circuit - Stimulus for EIS
V_source 100 0 AC 1V
X_cell 100 0 RandlesCell

* AC Analysis settings
.ac dec 10 0.001 10000000000.0

.control
  run
  set units = si
  
  * Define the Frequency vector
  let freq = frequency
  
  * Calculate Complex Impedance
  * Note: I(V_source) is negative convention in SPICE, so we use -I to get positive Z
  let Z = V(100) / -I(V_source)
  
  * Extract Components for EIS Analysis
  let Z_mag = abs(Z)
  let Z_phase = ph(Z)
  let Z_real = real(Z)
  let Z_imag = imag(Z)
  
  * Output to console (for parsing)
  print freq Z_mag Z_phase
  
  * Save data to file
  wrdata eis_data.txt Z_real Z_imag Z_mag Z_phase

.endc

.end
